module equals(output reg [55:0] out, input [55:0] in);
    initial begin
        assign out = in;
    end
endmodule



