module enot(output reg e_o, input e);
    initial begin
        assign e_o = ~e;
    end
endmodule



