module expansion(input [31:0] in, output [47:0] out);
    assign out = 48'b1;
endmodule
