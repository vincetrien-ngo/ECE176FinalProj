module equals #(parameter N=56)(output [N-1:0] out, input [N-1:0] in);


assign out = in;
endmodule




