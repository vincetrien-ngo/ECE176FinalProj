module equals(output reg [63:0] out, input [63:0] in);
    initial begin
        assign out = in;
    end
endmodule



