module equals_kb_ks(output reg [55:0] kp, input [55:0] ks);
    initial begin
        assign kp = ks;
    end
endmodule


