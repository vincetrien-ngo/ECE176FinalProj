
module main();

endmodule
