module equals(out, in);
parameter N=56;
output [N-1:0] out;
inout [N-1:0] in;
assign out = in;
endmodule




